`timescale 1ns / 1ps

module testbench;

    //arbiter_test arbiter_test();
    //testA test_A();
    testB test_B();
    //testC test_C();
    testC8 test_C8();

endmodule